Testje


V1 1 0 DC 8
R1 1 2 2
R2 2 0 4
I1 2 3 1
R3 3 4 6
V2 0 4 5
R4 3 5 9
R5 5 4 15
*VMEAS 5 4 0

.op
.end
